`timescale 1us/1ns

module tb_mux_4x_nbit();

	parameter BUS_WIDTH = 8;
	reg [BUS_WIDTH-1:0] a;
	reg [BUS_WIDTH-1:0] b;
	reg [BUS_WIDTH-1:0] c;
	reg [BUS_WIDTH-1:0] d;
	reg [1:0] sel;
	wire [BUS_WIDTH-1:0] y;
	
	integer i;

	// Instantiate the DUT
	mux_4x_nbit #(.BUS_WIDTH(BUS_WIDTH)) MUX0 (
		.a(a),
		.b(b),
		.c(c),
		.d(d),
		.sel(sel),
		.y(y)
	);

	initial begin
		$monitor($time, " a = %0d, b = %0d, c = %0d, d = %0d, sel = %0d, y = %0d", a, b, c, d, sel, y);

		#1; sel = 0; a = 0; b = 0;  c = 0; d = 0;

		for (i = 0; i < 8; i = i + 1) begin
			#1;
			sel = $urandom() % 4;
			a = $urandom() % 256;
			b = $urandom() % 256;
			c = $urandom() % 256;
			d = $urandom() % 256;
		end
	end
endmodule
