module demux_nbit_x4
